`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   10:12:37 03/05/2019
// Design Name:   traffic_light_controller
// Module Name:   Z:/shared_folder/cs141/pa3/lab3_start/test_traffic_light_controller.v
// Project Name:  lab3_start
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: traffic_light_controller
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test_traffic_light_controller;

	// Inputs
	reg clk;
	reg rst;
	wire [3:0] timer_out; // originally reg.
	reg car_ns;
	reg car_ew;
	reg ped;

	// Outputs
	wire timer_en;
	wire timer_load;
	wire [3:0] timer_init;
	wire [2:0] light_ns;
	wire [2:0] light_ew;
	wire [1:0] light_ped;
	
	// clk is 1 second clock generated by the testbench

	// Instantiate Timer 
	timer timer (
		.clk(clk),
		.rst(rst),
		.en(timer_en),
		.load(timer_load),
		.init(timer_init),
		.out(timer_out)
	);

	// Instantiate the Unit Under Test (UUT)
	traffic_light_controller uut (
		.clk(clk), 
		.rst(rst), 
		.timer_en(timer_en), 
		.timer_load(timer_load), 
		.timer_init(timer_init), 
		.timer_out(timer_out), 
		.car_ns(car_ns), 
		.car_ew(car_ew), 
		.ped(ped), 
		.light_ns(light_ns), 
		.light_ew(light_ew), 
		.light_ped(light_ped)
	);

	integer timepassed = 4'd0;
	integer T = 32'd1000000000; // 1 second period
	integer i;
	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 0;
		car_ns = 0;
		car_ew = 0;
		ped = 0;

		//Wait a bit and reset
		for(i = 0; i < 5; i = i + 1) begin
			#(T);
		end
		rst = 1;
		#T;
		rst = 0;
		
		for(i = 0; i < 24; i = i + 1) begin
			#(T);
		end
      
		ped = !ped;	//pedestrian arrives
		
		for(i = 0; i < 20; i = i + 1) begin
			#(T);
		end
		
		ped = !ped;	//ped leaves
		car_ns = !car_ns;	//cars arrive on both
		car_ew = !car_ew;

		for(i = 0; i < 10; i = i + 1) begin
			#(T);
		end
		
		car_ew = !car_ew;	//cars leave ew
		
		for(i = 0; i < 20; i = i + 1) begin
			#(T);
		end
		
		car_ns = !car_ns;	//cars leave ns
		
		for(i = 0; i < 20; i = i + 1) begin
			#(T);
		end
		
		$finish;

	end
	
	reg[7:0] cur;
	reg[7:0] prev;
	
	//Run a clock

	always begin
		#(T/2);
		clk = 1'b0;
		#(T/2);
		clk = 1'b1;
		timepassed = timepassed + 1;
	end
	
	// Test blocks checking requirements
	always @(light_ns, light_ew, light_ped) begin
		#2;
		prev = cur;
		cur = {light_ns, light_ped, light_ew};
	
		
		$display("TIME = %d	STATE = %b", timepassed, cur[7:0]);
		case(prev)
			8'b00100001 : begin	//test for transition to ped
				if(cur[7:0] !== 8'b00111001) begin
					$display("ERROR: Rule 2  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
			end
			8'b00111001 : begin	//test for transition to green light
				if(cur[7:0] == 8'b00100001) begin
					$display("Warning: Reset  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
				else if(cur[7:0] !== 8'b10010001 && cur[7:0] !== 8'b00101100) begin
					$display("%b", cur[7:0]);
					$display("Warning: Rule 4 (not lights)  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
				if(car_ns == 1 && cur[7:0] !== 8'b10010001) begin
					$display("Warning: Rule 4 (car waiting NS)  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
				if(car_ew == 1 && cur[7:0] !== 8'b00101100) begin
					$display("Warning: Rule 4 (car waiting EW)  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
			end

			8'b10010001: begin	// test for transition to yellow
				if(cur[7:0] !== 8'b01010001) begin
					$display("ERROR: Rule 8 (NS)  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
			end
			
			8'b00101100: begin	// test for transition to yellow
				if(cur !== 8'b00101010) begin
					$display("ERROR: Rule 8 (NS)  Cur: NS=%b, EW=%b, PED=%b		Prev: NS=%b, EW=%b, PED=%b		Time=%b", cur[7:5], cur[2:0], cur[4:3], prev[7:5], prev[2:0], prev[4:3], timepassed);
				end
			end
			
		endcase		
		
	end
      
endmodule

